//and gate coding
//added extra line after clone to do pull in local repo

module and_g(y,a,b);
	input a,b;
	output wire y;

	assign y=a&b;


endmodule
