//and gate coding

module and_g(y,a,b);
	input a,b;
	output wire y;

	assign y=a&b;


endmodule
